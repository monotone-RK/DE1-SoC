/******************************************************************************/
/* Clock & Reset Generator                                                    */
/******************************************************************************/

`default_nettype none

/* Clock Generator                                                            */
/******************************************************************************/
module clockgen(// interface 'refclk'
	        input wire refclk,
	        // interface 'reset'
	        input wire rst,
                
	        // interface 'outclk0'
	        output wire outclk_0,
	        // interface 'locked'
	        output wire locked);
  
  altera_pll #(
	       .fractional_vco_multiplier("false"),
	       .reference_clock_frequency("50.0 MHz"),
	       .operation_mode("normal"),
	       .number_of_clocks(1),
	       .output_clock_frequency0("100.000000 MHz"),
	       .phase_shift0("0 ps"),
	       .duty_cycle0(50),
	       .output_clock_frequency1("0 MHz"),
	       .phase_shift1("0 ps"),
	       .duty_cycle1(50),
	       .output_clock_frequency2("0 MHz"),
	       .phase_shift2("0 ps"),
	       .duty_cycle2(50),
	       .output_clock_frequency3("0 MHz"),
	       .phase_shift3("0 ps"),
	       .duty_cycle3(50),
	       .output_clock_frequency4("0 MHz"),
	       .phase_shift4("0 ps"),
	       .duty_cycle4(50),
	       .output_clock_frequency5("0 MHz"),
	       .phase_shift5("0 ps"),
	       .duty_cycle5(50),
	       .output_clock_frequency6("0 MHz"),
	       .phase_shift6("0 ps"),
	       .duty_cycle6(50),
	       .output_clock_frequency7("0 MHz"),
	       .phase_shift7("0 ps"),
	       .duty_cycle7(50),
	       .output_clock_frequency8("0 MHz"),
	       .phase_shift8("0 ps"),
	       .duty_cycle8(50),
	       .output_clock_frequency9("0 MHz"),
	       .phase_shift9("0 ps"),
	       .duty_cycle9(50),
	       .output_clock_frequency10("0 MHz"),
	       .phase_shift10("0 ps"),
	       .duty_cycle10(50),
	       .output_clock_frequency11("0 MHz"),
	       .phase_shift11("0 ps"),
	       .duty_cycle11(50),
	       .output_clock_frequency12("0 MHz"),
	       .phase_shift12("0 ps"),
	       .duty_cycle12(50),
	       .output_clock_frequency13("0 MHz"),
	       .phase_shift13("0 ps"),
	       .duty_cycle13(50),
	       .output_clock_frequency14("0 MHz"),
	       .phase_shift14("0 ps"),
	       .duty_cycle14(50),
	       .output_clock_frequency15("0 MHz"),
	       .phase_shift15("0 ps"),
	       .duty_cycle15(50),
	       .output_clock_frequency16("0 MHz"),
	       .phase_shift16("0 ps"),
	       .duty_cycle16(50),
	       .output_clock_frequency17("0 MHz"),
	       .phase_shift17("0 ps"),
	       .duty_cycle17(50),
	       .pll_type("General"),
	       .pll_subtype("General")
	       ) 
  altera_pll_i (
		.rst	(rst),
		.outclk	({outclk_0}),
		.locked	(locked),
		.fboutclk	( ),
		.fbclk	(1'b0),
		.refclk	(refclk)
	        );
endmodule

/* Reset Generator :  generate about 100 cycle reset signal                   */
/******************************************************************************/
module resetgen(input  wire CLK, 
                input  wire RST_X_I, 
                output wire RST_X_O);

  reg [7:0] cnt;
  assign RST_X_O = cnt[7];

  always @(posedge CLK) begin
    if      (!RST_X_I) cnt <= 0;
    else if (~RST_X_O) cnt <= (cnt + 1'b1);
  end
endmodule

/******************************************************************************/
module CLKRSTGEN(input  wire CLK_I, 
                 input  wire RST_X_I, 
                 output wire CLK_O, 
                 output wire RST_X_O);

  wire LOCKED;
  clockgen clkgen(.refclk(CLK_I),
                  .rst(~RST_X_I),
                  .outclk_0(CLK_O), 
                  .locked(LOCKED));
  resetgen rstgen(CLK_O, LOCKED, RST_X_O);
endmodule

`default_nettype wire
